`define DATA_WIDTH 8
`define CMD_WIDTH 4
`define N $clog2(`DATA_WIDTH)
`define no_of_trans 500
